// fpga_sdram_controller.v

// Generated using ACDS version 13.0sp1 232 at 2015.08.08.23:10:11

`timescale 1 ps / 1 ps
module fpga_sdram_controller (
		input  wire        clk_clk,                      //                  clk.clk
		input  wire        reset_reset_n,                //                reset.reset_n
		output wire [12:0] memory_mem_a,                 //               memory.mem_a
		output wire [2:0]  memory_mem_ba,                //                     .mem_ba
		output wire [0:0]  memory_mem_ck,                //                     .mem_ck
		output wire [0:0]  memory_mem_ck_n,              //                     .mem_ck_n
		output wire [0:0]  memory_mem_cke,               //                     .mem_cke
		output wire [0:0]  memory_mem_cs_n,              //                     .mem_cs_n
		output wire [3:0]  memory_mem_dm,                //                     .mem_dm
		output wire [0:0]  memory_mem_ras_n,             //                     .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,             //                     .mem_cas_n
		output wire [0:0]  memory_mem_we_n,              //                     .mem_we_n
		output wire        memory_mem_reset_n,           //                     .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                //                     .mem_dq
		inout  wire [3:0]  memory_mem_dqs,               //                     .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,             //                     .mem_dqs_n
		output wire [0:0]  memory_mem_odt,               //                     .mem_odt
		input  wire        oct_rzqin,                    //                  oct.rzqin
		input  wire [3:0]  axi_translator_slave_awid,    // axi_translator_slave.awid
		input  wire [31:0] axi_translator_slave_awaddr,  //                     .awaddr
		input  wire [7:0]  axi_translator_slave_awlen,   //                     .awlen
		input  wire [2:0]  axi_translator_slave_awsize,  //                     .awsize
		input  wire [1:0]  axi_translator_slave_awburst, //                     .awburst
		input  wire [0:0]  axi_translator_slave_awlock,  //                     .awlock
		input  wire [3:0]  axi_translator_slave_awcache, //                     .awcache
		input  wire [2:0]  axi_translator_slave_awprot,  //                     .awprot
		input  wire        axi_translator_slave_awvalid, //                     .awvalid
		output wire        axi_translator_slave_awready, //                     .awready
		input  wire [31:0] axi_translator_slave_wdata,   //                     .wdata
		input  wire [3:0]  axi_translator_slave_wstrb,   //                     .wstrb
		input  wire        axi_translator_slave_wlast,   //                     .wlast
		input  wire        axi_translator_slave_wvalid,  //                     .wvalid
		output wire        axi_translator_slave_wready,  //                     .wready
		output wire [3:0]  axi_translator_slave_bid,     //                     .bid
		output wire [1:0]  axi_translator_slave_bresp,   //                     .bresp
		output wire        axi_translator_slave_bvalid,  //                     .bvalid
		input  wire        axi_translator_slave_bready,  //                     .bready
		input  wire [3:0]  axi_translator_slave_arid,    //                     .arid
		input  wire [31:0] axi_translator_slave_araddr,  //                     .araddr
		input  wire [7:0]  axi_translator_slave_arlen,   //                     .arlen
		input  wire [2:0]  axi_translator_slave_arsize,  //                     .arsize
		input  wire [1:0]  axi_translator_slave_arburst, //                     .arburst
		input  wire [0:0]  axi_translator_slave_arlock,  //                     .arlock
		input  wire [3:0]  axi_translator_slave_arcache, //                     .arcache
		input  wire [2:0]  axi_translator_slave_arprot,  //                     .arprot
		input  wire        axi_translator_slave_arvalid, //                     .arvalid
		output wire        axi_translator_slave_arready, //                     .arready
		output wire [3:0]  axi_translator_slave_rid,     //                     .rid
		output wire [31:0] axi_translator_slave_rdata,   //                     .rdata
		output wire [1:0]  axi_translator_slave_rresp,   //                     .rresp
		output wire        axi_translator_slave_rlast,   //                     .rlast
		output wire        axi_translator_slave_rvalid,  //                     .rvalid
		input  wire        axi_translator_slave_rready   //                     .rready
	);

	wire          axi_translator_m0_awvalid;                                                                   // axi_translator:m0_awvalid -> axi_translator_m0_translator:s0_awvalid
	wire    [2:0] axi_translator_m0_arsize;                                                                    // axi_translator:m0_arsize -> axi_translator_m0_translator:s0_arsize
	wire    [0:0] axi_translator_m0_arlock;                                                                    // axi_translator:m0_arlock -> axi_translator_m0_translator:s0_arlock
	wire    [3:0] axi_translator_m0_awcache;                                                                   // axi_translator:m0_awcache -> axi_translator_m0_translator:s0_awcache
	wire          axi_translator_m0_arready;                                                                   // axi_translator_m0_translator:s0_arready -> axi_translator:m0_arready
	wire    [3:0] axi_translator_m0_arqos;                                                                     // axi_translator:m0_arqos -> axi_translator_m0_translator:s0_arqos
	wire    [7:0] axi_translator_m0_arid;                                                                      // axi_translator:m0_arid -> axi_translator_m0_translator:s0_arid
	wire          axi_translator_m0_rready;                                                                    // axi_translator:m0_rready -> axi_translator_m0_translator:s0_rready
	wire    [3:0] axi_translator_m0_arregion;                                                                  // axi_translator:m0_arregion -> axi_translator_m0_translator:s0_arregion
	wire          axi_translator_m0_bready;                                                                    // axi_translator:m0_bready -> axi_translator_m0_translator:s0_bready
	wire    [2:0] axi_translator_m0_awsize;                                                                    // axi_translator:m0_awsize -> axi_translator_m0_translator:s0_awsize
	wire    [2:0] axi_translator_m0_awprot;                                                                    // axi_translator:m0_awprot -> axi_translator_m0_translator:s0_awprot
	wire          axi_translator_m0_arvalid;                                                                   // axi_translator:m0_arvalid -> axi_translator_m0_translator:s0_arvalid
	wire    [3:0] axi_translator_m0_awqos;                                                                     // axi_translator:m0_awqos -> axi_translator_m0_translator:s0_awqos
	wire    [2:0] axi_translator_m0_arprot;                                                                    // axi_translator:m0_arprot -> axi_translator_m0_translator:s0_arprot
	wire    [7:0] axi_translator_m0_bid;                                                                       // axi_translator_m0_translator:s0_bid -> axi_translator:m0_bid
	wire    [7:0] axi_translator_m0_arlen;                                                                     // axi_translator:m0_arlen -> axi_translator_m0_translator:s0_arlen
	wire          axi_translator_m0_awready;                                                                   // axi_translator_m0_translator:s0_awready -> axi_translator:m0_awready
	wire    [7:0] axi_translator_m0_awid;                                                                      // axi_translator:m0_awid -> axi_translator_m0_translator:s0_awid
	wire          axi_translator_m0_bvalid;                                                                    // axi_translator_m0_translator:s0_bvalid -> axi_translator:m0_bvalid
	wire    [3:0] axi_translator_m0_awregion;                                                                  // axi_translator:m0_awregion -> axi_translator_m0_translator:s0_awregion
	wire    [0:0] axi_translator_m0_awlock;                                                                    // axi_translator:m0_awlock -> axi_translator_m0_translator:s0_awlock
	wire    [1:0] axi_translator_m0_awburst;                                                                   // axi_translator:m0_awburst -> axi_translator_m0_translator:s0_awburst
	wire    [1:0] axi_translator_m0_bresp;                                                                     // axi_translator_m0_translator:s0_bresp -> axi_translator:m0_bresp
	wire    [3:0] axi_translator_m0_wstrb;                                                                     // axi_translator:m0_wstrb -> axi_translator_m0_translator:s0_wstrb
	wire          axi_translator_m0_rvalid;                                                                    // axi_translator_m0_translator:s0_rvalid -> axi_translator:m0_rvalid
	wire    [1:0] axi_translator_m0_arburst;                                                                   // axi_translator:m0_arburst -> axi_translator_m0_translator:s0_arburst
	wire   [31:0] axi_translator_m0_wdata;                                                                     // axi_translator:m0_wdata -> axi_translator_m0_translator:s0_wdata
	wire          axi_translator_m0_wready;                                                                    // axi_translator_m0_translator:s0_wready -> axi_translator:m0_wready
	wire   [31:0] axi_translator_m0_rdata;                                                                     // axi_translator_m0_translator:s0_rdata -> axi_translator:m0_rdata
	wire   [31:0] axi_translator_m0_araddr;                                                                    // axi_translator:m0_araddr -> axi_translator_m0_translator:s0_araddr
	wire    [3:0] axi_translator_m0_arcache;                                                                   // axi_translator:m0_arcache -> axi_translator_m0_translator:s0_arcache
	wire    [7:0] axi_translator_m0_awlen;                                                                     // axi_translator:m0_awlen -> axi_translator_m0_translator:s0_awlen
	wire   [31:0] axi_translator_m0_awaddr;                                                                    // axi_translator:m0_awaddr -> axi_translator_m0_translator:s0_awaddr
	wire    [7:0] axi_translator_m0_rid;                                                                       // axi_translator_m0_translator:s0_rid -> axi_translator:m0_rid
	wire          axi_translator_m0_wvalid;                                                                    // axi_translator:m0_wvalid -> axi_translator_m0_translator:s0_wvalid
	wire    [1:0] axi_translator_m0_rresp;                                                                     // axi_translator_m0_translator:s0_rresp -> axi_translator:m0_rresp
	wire          axi_translator_m0_wlast;                                                                     // axi_translator:m0_wlast -> axi_translator_m0_translator:s0_wlast
	wire          axi_translator_m0_rlast;                                                                     // axi_translator_m0_translator:s0_rlast -> axi_translator:m0_rlast
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_waitrequest;                           // mem_if_ddr3_emif_0:avl_ready -> mem_if_ddr3_emif_0_avl_translator:av_waitrequest
	wire    [5:0] mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_burstcount;                            // mem_if_ddr3_emif_0_avl_translator:av_burstcount -> mem_if_ddr3_emif_0:avl_size
	wire  [127:0] mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_writedata;                             // mem_if_ddr3_emif_0_avl_translator:av_writedata -> mem_if_ddr3_emif_0:avl_wdata
	wire   [23:0] mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_address;                               // mem_if_ddr3_emif_0_avl_translator:av_address -> mem_if_ddr3_emif_0:avl_addr
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_write;                                 // mem_if_ddr3_emif_0_avl_translator:av_write -> mem_if_ddr3_emif_0:avl_write_req
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_beginbursttransfer;                    // mem_if_ddr3_emif_0_avl_translator:av_beginbursttransfer -> mem_if_ddr3_emif_0:avl_burstbegin
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_read;                                  // mem_if_ddr3_emif_0_avl_translator:av_read -> mem_if_ddr3_emif_0:avl_read_req
	wire  [127:0] mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_readdata;                              // mem_if_ddr3_emif_0:avl_rdata -> mem_if_ddr3_emif_0_avl_translator:av_readdata
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_readdatavalid;                         // mem_if_ddr3_emif_0:avl_rdata_valid -> mem_if_ddr3_emif_0_avl_translator:av_readdatavalid
	wire   [15:0] mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_byteenable;                            // mem_if_ddr3_emif_0_avl_translator:av_byteenable -> mem_if_ddr3_emif_0:avl_be
	wire          mem_if_ddr3_emif_0_afi_clk_clk;                                                              // mem_if_ddr3_emif_0:afi_clk -> [burst_adapter:clk, cmd_xbar_mux:clk, crosser:out_clk, crosser_001:out_clk, crosser_002:in_clk, crosser_003:in_clk, id_router:clk, mem_if_ddr3_emif_0_avl_translator:clk, mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:clk, mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rst_controller_001:clk, width_adapter:clk]
	wire          axi_translator_m0_translator_m0_awvalid;                                                     // axi_translator_m0_translator:m0_awvalid -> axi_translator_m0_translator_m0_agent:awvalid
	wire    [2:0] axi_translator_m0_translator_m0_arsize;                                                      // axi_translator_m0_translator:m0_arsize -> axi_translator_m0_translator_m0_agent:arsize
	wire    [0:0] axi_translator_m0_translator_m0_buser;                                                       // axi_translator_m0_translator_m0_agent:buser -> axi_translator_m0_translator:m0_buser
	wire    [0:0] axi_translator_m0_translator_m0_arlock;                                                      // axi_translator_m0_translator:m0_arlock -> axi_translator_m0_translator_m0_agent:arlock
	wire    [3:0] axi_translator_m0_translator_m0_awcache;                                                     // axi_translator_m0_translator:m0_awcache -> axi_translator_m0_translator_m0_agent:awcache
	wire          axi_translator_m0_translator_m0_arready;                                                     // axi_translator_m0_translator_m0_agent:arready -> axi_translator_m0_translator:m0_arready
	wire    [3:0] axi_translator_m0_translator_m0_arqos;                                                       // axi_translator_m0_translator:m0_arqos -> axi_translator_m0_translator_m0_agent:arqos
	wire    [7:0] axi_translator_m0_translator_m0_arid;                                                        // axi_translator_m0_translator:m0_arid -> axi_translator_m0_translator_m0_agent:arid
	wire          axi_translator_m0_translator_m0_rready;                                                      // axi_translator_m0_translator:m0_rready -> axi_translator_m0_translator_m0_agent:rready
	wire    [3:0] axi_translator_m0_translator_m0_arregion;                                                    // axi_translator_m0_translator:m0_arregion -> axi_translator_m0_translator_m0_agent:arregion
	wire    [0:0] axi_translator_m0_translator_m0_ruser;                                                       // axi_translator_m0_translator_m0_agent:ruser -> axi_translator_m0_translator:m0_ruser
	wire          axi_translator_m0_translator_m0_bready;                                                      // axi_translator_m0_translator:m0_bready -> axi_translator_m0_translator_m0_agent:bready
	wire    [2:0] axi_translator_m0_translator_m0_awsize;                                                      // axi_translator_m0_translator:m0_awsize -> axi_translator_m0_translator_m0_agent:awsize
	wire    [2:0] axi_translator_m0_translator_m0_awprot;                                                      // axi_translator_m0_translator:m0_awprot -> axi_translator_m0_translator_m0_agent:awprot
	wire          axi_translator_m0_translator_m0_arvalid;                                                     // axi_translator_m0_translator:m0_arvalid -> axi_translator_m0_translator_m0_agent:arvalid
	wire    [3:0] axi_translator_m0_translator_m0_awqos;                                                       // axi_translator_m0_translator:m0_awqos -> axi_translator_m0_translator_m0_agent:awqos
	wire    [2:0] axi_translator_m0_translator_m0_arprot;                                                      // axi_translator_m0_translator:m0_arprot -> axi_translator_m0_translator_m0_agent:arprot
	wire    [7:0] axi_translator_m0_translator_m0_arlen;                                                       // axi_translator_m0_translator:m0_arlen -> axi_translator_m0_translator_m0_agent:arlen
	wire    [7:0] axi_translator_m0_translator_m0_bid;                                                         // axi_translator_m0_translator_m0_agent:bid -> axi_translator_m0_translator:m0_bid
	wire          axi_translator_m0_translator_m0_awready;                                                     // axi_translator_m0_translator_m0_agent:awready -> axi_translator_m0_translator:m0_awready
	wire    [7:0] axi_translator_m0_translator_m0_awid;                                                        // axi_translator_m0_translator:m0_awid -> axi_translator_m0_translator_m0_agent:awid
	wire          axi_translator_m0_translator_m0_bvalid;                                                      // axi_translator_m0_translator_m0_agent:bvalid -> axi_translator_m0_translator:m0_bvalid
	wire    [3:0] axi_translator_m0_translator_m0_awregion;                                                    // axi_translator_m0_translator:m0_awregion -> axi_translator_m0_translator_m0_agent:awregion
	wire    [0:0] axi_translator_m0_translator_m0_awlock;                                                      // axi_translator_m0_translator:m0_awlock -> axi_translator_m0_translator_m0_agent:awlock
	wire    [1:0] axi_translator_m0_translator_m0_awburst;                                                     // axi_translator_m0_translator:m0_awburst -> axi_translator_m0_translator_m0_agent:awburst
	wire    [1:0] axi_translator_m0_translator_m0_bresp;                                                       // axi_translator_m0_translator_m0_agent:bresp -> axi_translator_m0_translator:m0_bresp
	wire    [0:0] axi_translator_m0_translator_m0_aruser;                                                      // axi_translator_m0_translator:m0_aruser -> axi_translator_m0_translator_m0_agent:aruser
	wire    [0:0] axi_translator_m0_translator_m0_awuser;                                                      // axi_translator_m0_translator:m0_awuser -> axi_translator_m0_translator_m0_agent:awuser
	wire    [3:0] axi_translator_m0_translator_m0_wstrb;                                                       // axi_translator_m0_translator:m0_wstrb -> axi_translator_m0_translator_m0_agent:wstrb
	wire          axi_translator_m0_translator_m0_rvalid;                                                      // axi_translator_m0_translator_m0_agent:rvalid -> axi_translator_m0_translator:m0_rvalid
	wire    [1:0] axi_translator_m0_translator_m0_arburst;                                                     // axi_translator_m0_translator:m0_arburst -> axi_translator_m0_translator_m0_agent:arburst
	wire   [31:0] axi_translator_m0_translator_m0_wdata;                                                       // axi_translator_m0_translator:m0_wdata -> axi_translator_m0_translator_m0_agent:wdata
	wire          axi_translator_m0_translator_m0_wready;                                                      // axi_translator_m0_translator_m0_agent:wready -> axi_translator_m0_translator:m0_wready
	wire   [31:0] axi_translator_m0_translator_m0_rdata;                                                       // axi_translator_m0_translator_m0_agent:rdata -> axi_translator_m0_translator:m0_rdata
	wire   [31:0] axi_translator_m0_translator_m0_araddr;                                                      // axi_translator_m0_translator:m0_araddr -> axi_translator_m0_translator_m0_agent:araddr
	wire    [3:0] axi_translator_m0_translator_m0_arcache;                                                     // axi_translator_m0_translator:m0_arcache -> axi_translator_m0_translator_m0_agent:arcache
	wire    [7:0] axi_translator_m0_translator_m0_awlen;                                                       // axi_translator_m0_translator:m0_awlen -> axi_translator_m0_translator_m0_agent:awlen
	wire   [31:0] axi_translator_m0_translator_m0_awaddr;                                                      // axi_translator_m0_translator:m0_awaddr -> axi_translator_m0_translator_m0_agent:awaddr
	wire    [0:0] axi_translator_m0_translator_m0_wuser;                                                       // axi_translator_m0_translator:m0_wuser -> axi_translator_m0_translator_m0_agent:wuser
	wire    [7:0] axi_translator_m0_translator_m0_rid;                                                         // axi_translator_m0_translator_m0_agent:rid -> axi_translator_m0_translator:m0_rid
	wire          axi_translator_m0_translator_m0_wvalid;                                                      // axi_translator_m0_translator:m0_wvalid -> axi_translator_m0_translator_m0_agent:wvalid
	wire    [1:0] axi_translator_m0_translator_m0_rresp;                                                       // axi_translator_m0_translator_m0_agent:rresp -> axi_translator_m0_translator:m0_rresp
	wire          axi_translator_m0_translator_m0_wlast;                                                       // axi_translator_m0_translator:m0_wlast -> axi_translator_m0_translator_m0_agent:wlast
	wire          axi_translator_m0_translator_m0_rlast;                                                       // axi_translator_m0_translator_m0_agent:rlast -> axi_translator_m0_translator:m0_rlast
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // mem_if_ddr3_emif_0_avl_translator:uav_waitrequest -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [9:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_burstcount -> mem_if_ddr3_emif_0_avl_translator:uav_burstcount
	wire  [127:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_writedata;               // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_writedata -> mem_if_ddr3_emif_0_avl_translator:uav_writedata
	wire   [31:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_address;                 // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_address -> mem_if_ddr3_emif_0_avl_translator:uav_address
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_write;                   // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_write -> mem_if_ddr3_emif_0_avl_translator:uav_write
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_lock;                    // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_lock -> mem_if_ddr3_emif_0_avl_translator:uav_lock
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_read;                    // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_read -> mem_if_ddr3_emif_0_avl_translator:uav_read
	wire  [127:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdata;                // mem_if_ddr3_emif_0_avl_translator:uav_readdata -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // mem_if_ddr3_emif_0_avl_translator:uav_readdatavalid -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mem_if_ddr3_emif_0_avl_translator:uav_debugaccess
	wire   [15:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:m0_byteenable -> mem_if_ddr3_emif_0_avl_translator:uav_byteenable
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_valid -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [233:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_data;             // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_data -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [233:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [129:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;       // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [129:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;        // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;       // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          axi_translator_m0_translator_m0_agent_write_cp_endofpacket;                                  // axi_translator_m0_translator_m0_agent:write_cp_endofpacket -> addr_router:sink_endofpacket
	wire          axi_translator_m0_translator_m0_agent_write_cp_valid;                                        // axi_translator_m0_translator_m0_agent:write_cp_valid -> addr_router:sink_valid
	wire          axi_translator_m0_translator_m0_agent_write_cp_startofpacket;                                // axi_translator_m0_translator_m0_agent:write_cp_startofpacket -> addr_router:sink_startofpacket
	wire  [124:0] axi_translator_m0_translator_m0_agent_write_cp_data;                                         // axi_translator_m0_translator_m0_agent:write_cp_data -> addr_router:sink_data
	wire          axi_translator_m0_translator_m0_agent_write_cp_ready;                                        // addr_router:sink_ready -> axi_translator_m0_translator_m0_agent:write_cp_ready
	wire          axi_translator_m0_translator_m0_agent_read_cp_endofpacket;                                   // axi_translator_m0_translator_m0_agent:read_cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          axi_translator_m0_translator_m0_agent_read_cp_valid;                                         // axi_translator_m0_translator_m0_agent:read_cp_valid -> addr_router_001:sink_valid
	wire          axi_translator_m0_translator_m0_agent_read_cp_startofpacket;                                 // axi_translator_m0_translator_m0_agent:read_cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [124:0] axi_translator_m0_translator_m0_agent_read_cp_data;                                          // axi_translator_m0_translator_m0_agent:read_cp_data -> addr_router_001:sink_data
	wire          axi_translator_m0_translator_m0_agent_read_cp_ready;                                         // addr_router_001:sink_ready -> axi_translator_m0_translator_m0_agent:read_cp_ready
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_valid;                   // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [232:0] mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_data;                    // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:rp_ready
	wire          burst_adapter_source0_endofpacket;                                                           // burst_adapter:source0_endofpacket -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                 // burst_adapter:source0_valid -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                         // burst_adapter:source0_startofpacket -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [232:0] burst_adapter_source0_data;                                                                  // burst_adapter:source0_data -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                 // mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire    [1:0] burst_adapter_source0_channel;                                                               // burst_adapter:source0_channel -> mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:cp_channel
	wire          width_adapter_cmd_source_endofpacket;                                                        // width_adapter:cmd_out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_cmd_source_valid;                                                              // width_adapter:cmd_out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_cmd_source_startofpacket;                                                      // width_adapter:cmd_out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [232:0] width_adapter_cmd_source_data;                                                               // width_adapter:cmd_out_data -> burst_adapter:sink0_data
	wire    [1:0] width_adapter_cmd_source_channel;                                                            // width_adapter:cmd_out_channel -> burst_adapter:sink0_channel
	wire          width_adapter_cmd_source_ready;                                                              // burst_adapter:sink0_ready -> width_adapter:cmd_out_ready
	wire          id_router_src_endofpacket;                                                                   // id_router:src_endofpacket -> width_adapter:rsp_in_endofpacket
	wire          id_router_src_valid;                                                                         // id_router:src_valid -> width_adapter:rsp_in_valid
	wire          id_router_src_startofpacket;                                                                 // id_router:src_startofpacket -> width_adapter:rsp_in_startofpacket
	wire  [232:0] id_router_src_data;                                                                          // id_router:src_data -> width_adapter:rsp_in_data
	wire    [1:0] id_router_src_channel;                                                                       // id_router:src_channel -> width_adapter:rsp_in_channel
	wire          id_router_src_ready;                                                                         // width_adapter:rsp_in_ready -> id_router:src_ready
	wire          rst_controller_reset_out_reset;                                                              // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, axi_translator:aresetn, axi_translator_m0_translator:aresetn, axi_translator_m0_translator_m0_agent:aresetn, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:out_reset, crosser_003:out_reset]
	wire          rst_controller_001_reset_out_reset;                                                          // rst_controller_001:reset_out -> [burst_adapter:reset, cmd_xbar_mux:reset, crosser:out_reset, crosser_001:out_reset, crosser_002:in_reset, crosser_003:in_reset, id_router:reset, mem_if_ddr3_emif_0_avl_translator:reset, mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent:reset, mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, width_adapter:reset]
	wire          mem_if_ddr3_emif_0_afi_reset_reset;                                                          // mem_if_ddr3_emif_0:afi_reset_n -> rst_controller_001:reset_in0
	wire          addr_router_src_endofpacket;                                                                 // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                       // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                               // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [124:0] addr_router_src_data;                                                                        // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire    [1:0] addr_router_src_channel;                                                                     // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                       // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          crosser_002_out_ready;                                                                       // axi_translator_m0_translator_m0_agent:write_rp_ready -> crosser_002:out_ready
	wire          addr_router_001_src_endofpacket;                                                             // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                   // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                           // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [124:0] addr_router_001_src_data;                                                                    // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire    [1:0] addr_router_001_src_channel;                                                                 // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                   // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          crosser_003_out_ready;                                                                       // axi_translator_m0_translator_m0_agent:read_rp_ready -> crosser_003:out_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                // cmd_xbar_mux:src_endofpacket -> width_adapter:cmd_in_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                      // cmd_xbar_mux:src_valid -> width_adapter:cmd_in_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                              // cmd_xbar_mux:src_startofpacket -> width_adapter:cmd_in_startofpacket
	wire  [124:0] cmd_xbar_mux_src_data;                                                                       // cmd_xbar_mux:src_data -> width_adapter:cmd_in_data
	wire    [1:0] cmd_xbar_mux_src_channel;                                                                    // cmd_xbar_mux:src_channel -> width_adapter:cmd_in_channel
	wire          cmd_xbar_mux_src_ready;                                                                      // width_adapter:cmd_in_ready -> cmd_xbar_mux:src_ready
	wire          width_adapter_rsp_source_endofpacket;                                                        // width_adapter:rsp_out_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          width_adapter_rsp_source_valid;                                                              // width_adapter:rsp_out_valid -> rsp_xbar_demux:sink_valid
	wire          width_adapter_rsp_source_startofpacket;                                                      // width_adapter:rsp_out_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [124:0] width_adapter_rsp_source_data;                                                               // width_adapter:rsp_out_data -> rsp_xbar_demux:sink_data
	wire    [1:0] width_adapter_rsp_source_channel;                                                            // width_adapter:rsp_out_channel -> rsp_xbar_demux:sink_channel
	wire          width_adapter_rsp_source_ready;                                                              // rsp_xbar_demux:sink_ready -> width_adapter:rsp_out_ready
	wire          crosser_out_endofpacket;                                                                     // crosser:out_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          crosser_out_valid;                                                                           // crosser:out_valid -> cmd_xbar_mux:sink0_valid
	wire          crosser_out_startofpacket;                                                                   // crosser:out_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [124:0] crosser_out_data;                                                                            // crosser:out_data -> cmd_xbar_mux:sink0_data
	wire    [1:0] crosser_out_channel;                                                                         // crosser:out_channel -> cmd_xbar_mux:sink0_channel
	wire          crosser_out_ready;                                                                           // cmd_xbar_mux:sink0_ready -> crosser:out_ready
	wire          cmd_xbar_demux_src0_endofpacket;                                                             // cmd_xbar_demux:src0_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                   // cmd_xbar_demux:src0_valid -> crosser:in_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                           // cmd_xbar_demux:src0_startofpacket -> crosser:in_startofpacket
	wire  [124:0] cmd_xbar_demux_src0_data;                                                                    // cmd_xbar_demux:src0_data -> crosser:in_data
	wire    [1:0] cmd_xbar_demux_src0_channel;                                                                 // cmd_xbar_demux:src0_channel -> crosser:in_channel
	wire          cmd_xbar_demux_src0_ready;                                                                   // crosser:in_ready -> cmd_xbar_demux:src0_ready
	wire          crosser_001_out_endofpacket;                                                                 // crosser_001:out_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          crosser_001_out_valid;                                                                       // crosser_001:out_valid -> cmd_xbar_mux:sink1_valid
	wire          crosser_001_out_startofpacket;                                                               // crosser_001:out_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [124:0] crosser_001_out_data;                                                                        // crosser_001:out_data -> cmd_xbar_mux:sink1_data
	wire    [1:0] crosser_001_out_channel;                                                                     // crosser_001:out_channel -> cmd_xbar_mux:sink1_channel
	wire          crosser_001_out_ready;                                                                       // cmd_xbar_mux:sink1_ready -> crosser_001:out_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                         // cmd_xbar_demux_001:src0_endofpacket -> crosser_001:in_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                               // cmd_xbar_demux_001:src0_valid -> crosser_001:in_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                       // cmd_xbar_demux_001:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [124:0] cmd_xbar_demux_001_src0_data;                                                                // cmd_xbar_demux_001:src0_data -> crosser_001:in_data
	wire    [1:0] cmd_xbar_demux_001_src0_channel;                                                             // cmd_xbar_demux_001:src0_channel -> crosser_001:in_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                               // crosser_001:in_ready -> cmd_xbar_demux_001:src0_ready
	wire          crosser_002_out_endofpacket;                                                                 // crosser_002:out_endofpacket -> axi_translator_m0_translator_m0_agent:write_rp_endofpacket
	wire          crosser_002_out_valid;                                                                       // crosser_002:out_valid -> axi_translator_m0_translator_m0_agent:write_rp_valid
	wire          crosser_002_out_startofpacket;                                                               // crosser_002:out_startofpacket -> axi_translator_m0_translator_m0_agent:write_rp_startofpacket
	wire  [124:0] crosser_002_out_data;                                                                        // crosser_002:out_data -> axi_translator_m0_translator_m0_agent:write_rp_data
	wire    [1:0] crosser_002_out_channel;                                                                     // crosser_002:out_channel -> axi_translator_m0_translator_m0_agent:write_rp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                             // rsp_xbar_demux:src0_endofpacket -> crosser_002:in_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                   // rsp_xbar_demux:src0_valid -> crosser_002:in_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                           // rsp_xbar_demux:src0_startofpacket -> crosser_002:in_startofpacket
	wire  [124:0] rsp_xbar_demux_src0_data;                                                                    // rsp_xbar_demux:src0_data -> crosser_002:in_data
	wire    [1:0] rsp_xbar_demux_src0_channel;                                                                 // rsp_xbar_demux:src0_channel -> crosser_002:in_channel
	wire          rsp_xbar_demux_src0_ready;                                                                   // crosser_002:in_ready -> rsp_xbar_demux:src0_ready
	wire          crosser_003_out_endofpacket;                                                                 // crosser_003:out_endofpacket -> axi_translator_m0_translator_m0_agent:read_rp_endofpacket
	wire          crosser_003_out_valid;                                                                       // crosser_003:out_valid -> axi_translator_m0_translator_m0_agent:read_rp_valid
	wire          crosser_003_out_startofpacket;                                                               // crosser_003:out_startofpacket -> axi_translator_m0_translator_m0_agent:read_rp_startofpacket
	wire  [124:0] crosser_003_out_data;                                                                        // crosser_003:out_data -> axi_translator_m0_translator_m0_agent:read_rp_data
	wire    [1:0] crosser_003_out_channel;                                                                     // crosser_003:out_channel -> axi_translator_m0_translator_m0_agent:read_rp_channel
	wire          rsp_xbar_demux_src1_endofpacket;                                                             // rsp_xbar_demux:src1_endofpacket -> crosser_003:in_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                   // rsp_xbar_demux:src1_valid -> crosser_003:in_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                           // rsp_xbar_demux:src1_startofpacket -> crosser_003:in_startofpacket
	wire  [124:0] rsp_xbar_demux_src1_data;                                                                    // rsp_xbar_demux:src1_data -> crosser_003:in_data
	wire    [1:0] rsp_xbar_demux_src1_channel;                                                                 // rsp_xbar_demux:src1_channel -> crosser_003:in_channel
	wire          rsp_xbar_demux_src1_ready;                                                                   // crosser_003:in_ready -> rsp_xbar_demux:src1_ready

	fpga_sdram_controller_mem_if_ddr3_emif_0 mem_if_ddr3_emif_0 (
		.pll_ref_clk               (clk_clk),                                                                  //      pll_ref_clk.clk
		.global_reset_n            (reset_reset_n),                                                            //     global_reset.reset_n
		.soft_reset_n              (reset_reset_n),                                                            //       soft_reset.reset_n
		.afi_clk                   (mem_if_ddr3_emif_0_afi_clk_clk),                                           //          afi_clk.clk
		.afi_half_clk              (),                                                                         //     afi_half_clk.clk
		.afi_reset_n               (mem_if_ddr3_emif_0_afi_reset_reset),                                       //        afi_reset.reset_n
		.afi_reset_export_n        (),                                                                         // afi_reset_export.reset_n
		.mem_a                     (memory_mem_a),                                                             //           memory.mem_a
		.mem_ba                    (memory_mem_ba),                                                            //                 .mem_ba
		.mem_ck                    (memory_mem_ck),                                                            //                 .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                                                          //                 .mem_ck_n
		.mem_cke                   (memory_mem_cke),                                                           //                 .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                                                          //                 .mem_cs_n
		.mem_dm                    (memory_mem_dm),                                                            //                 .mem_dm
		.mem_ras_n                 (memory_mem_ras_n),                                                         //                 .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                                                         //                 .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                                                          //                 .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),                                                       //                 .mem_reset_n
		.mem_dq                    (memory_mem_dq),                                                            //                 .mem_dq
		.mem_dqs                   (memory_mem_dqs),                                                           //                 .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                                                         //                 .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                                                           //                 .mem_odt
		.avl_ready                 (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin            (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_address),            //                 .address
		.avl_rdata_valid           (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_readdata),           //                 .readdata
		.avl_wdata                 (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_writedata),          //                 .writedata
		.avl_be                    (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_byteenable),         //                 .byteenable
		.avl_read_req              (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_read),               //                 .read
		.avl_write_req             (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_write),              //                 .write
		.avl_size                  (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_burstcount),         //                 .burstcount
		.local_init_done           (),                                                                         //           status.local_init_done
		.local_cal_success         (),                                                                         //                 .local_cal_success
		.local_cal_fail            (),                                                                         //                 .local_cal_fail
		.oct_rzqin                 (oct_rzqin),                                                                //              oct.rzqin
		.pll_mem_clk               (),                                                                         //      pll_sharing.pll_mem_clk
		.pll_write_clk             (),                                                                         //                 .pll_write_clk
		.pll_write_clk_pre_phy_clk (),                                                                         //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (),                                                                         //                 .pll_addr_cmd_clk
		.pll_locked                (),                                                                         //                 .pll_locked
		.pll_avl_clk               (),                                                                         //                 .pll_avl_clk
		.pll_config_clk            (),                                                                         //                 .pll_config_clk
		.pll_mem_phy_clk           (),                                                                         //                 .pll_mem_phy_clk
		.afi_phy_clk               (),                                                                         //                 .afi_phy_clk
		.pll_avl_phy_clk           ()                                                                          //                 .pll_avl_phy_clk
	);

	altera_merlin_axi_translator #(
		.USE_S0_AWID                       (1),
		.USE_S0_AWREGION                   (0),
		.USE_M0_AWREGION                   (1),
		.USE_S0_AWLEN                      (1),
		.USE_S0_AWSIZE                     (1),
		.USE_S0_AWBURST                    (1),
		.USE_S0_AWLOCK                     (1),
		.USE_M0_AWLOCK                     (1),
		.USE_S0_AWCACHE                    (1),
		.USE_M0_AWCACHE                    (1),
		.USE_M0_AWPROT                     (1),
		.USE_S0_AWQOS                      (0),
		.USE_M0_AWQOS                      (1),
		.USE_S0_WSTRB                      (1),
		.USE_M0_WLAST                      (1),
		.USE_S0_BID                        (1),
		.USE_S0_BRESP                      (1),
		.USE_M0_BRESP                      (1),
		.USE_S0_ARID                       (1),
		.USE_S0_ARREGION                   (0),
		.USE_M0_ARREGION                   (1),
		.USE_S0_ARLEN                      (1),
		.USE_S0_ARSIZE                     (1),
		.USE_S0_ARBURST                    (1),
		.USE_S0_ARLOCK                     (1),
		.USE_M0_ARLOCK                     (1),
		.USE_M0_ARCACHE                    (1),
		.USE_M0_ARQOS                      (1),
		.USE_M0_ARPROT                     (1),
		.USE_S0_ARCACHE                    (1),
		.USE_S0_ARQOS                      (0),
		.USE_S0_RID                        (1),
		.USE_S0_RRESP                      (1),
		.USE_M0_RRESP                      (1),
		.USE_S0_RLAST                      (1),
		.M0_ID_WIDTH                       (8),
		.DATA_WIDTH                        (32),
		.S0_ID_WIDTH                       (4),
		.M0_ADDR_WIDTH                     (32),
		.S0_WRITE_ADDR_USER_WIDTH          (64),
		.S0_READ_ADDR_USER_WIDTH           (64),
		.M0_WRITE_ADDR_USER_WIDTH          (64),
		.M0_READ_ADDR_USER_WIDTH           (64),
		.S0_WRITE_DATA_USER_WIDTH          (64),
		.S0_WRITE_RESPONSE_DATA_USER_WIDTH (64),
		.S0_READ_DATA_USER_WIDTH           (64),
		.M0_WRITE_DATA_USER_WIDTH          (64),
		.M0_WRITE_RESPONSE_DATA_USER_WIDTH (64),
		.M0_READ_DATA_USER_WIDTH           (64),
		.S0_ADDR_WIDTH                     (32),
		.USE_S0_AWUSER                     (0),
		.USE_S0_ARUSER                     (0),
		.USE_S0_WUSER                      (0),
		.USE_S0_RUSER                      (0),
		.USE_S0_BUSER                      (0),
		.USE_M0_AWUSER                     (0),
		.USE_M0_ARUSER                     (0),
		.USE_M0_WUSER                      (0),
		.USE_M0_RUSER                      (0),
		.USE_M0_BUSER                      (0),
		.M0_AXI_VERSION                    ("AXI4"),
		.M0_BURST_LENGTH_WIDTH             (8),
		.S0_BURST_LENGTH_WIDTH             (8),
		.M0_LOCK_WIDTH                     (1),
		.S0_LOCK_WIDTH                     (1),
		.S0_AXI_VERSION                    ("AXI4")
	) axi_translator (
		.aclk        (clk_clk),                                                              //       clk.clk
		.aresetn     (~rst_controller_reset_out_reset),                                      // clk_reset.reset_n
		.s0_awid     (axi_translator_slave_awid),                                            //        s0.awid
		.s0_awaddr   (axi_translator_slave_awaddr),                                          //          .awaddr
		.s0_awlen    (axi_translator_slave_awlen),                                           //          .awlen
		.s0_awsize   (axi_translator_slave_awsize),                                          //          .awsize
		.s0_awburst  (axi_translator_slave_awburst),                                         //          .awburst
		.s0_awlock   (axi_translator_slave_awlock),                                          //          .awlock
		.s0_awcache  (axi_translator_slave_awcache),                                         //          .awcache
		.s0_awprot   (axi_translator_slave_awprot),                                          //          .awprot
		.s0_awvalid  (axi_translator_slave_awvalid),                                         //          .awvalid
		.s0_awready  (axi_translator_slave_awready),                                         //          .awready
		.s0_wdata    (axi_translator_slave_wdata),                                           //          .wdata
		.s0_wstrb    (axi_translator_slave_wstrb),                                           //          .wstrb
		.s0_wlast    (axi_translator_slave_wlast),                                           //          .wlast
		.s0_wvalid   (axi_translator_slave_wvalid),                                          //          .wvalid
		.s0_wready   (axi_translator_slave_wready),                                          //          .wready
		.s0_bid      (axi_translator_slave_bid),                                             //          .bid
		.s0_bresp    (axi_translator_slave_bresp),                                           //          .bresp
		.s0_bvalid   (axi_translator_slave_bvalid),                                          //          .bvalid
		.s0_bready   (axi_translator_slave_bready),                                          //          .bready
		.s0_arid     (axi_translator_slave_arid),                                            //          .arid
		.s0_araddr   (axi_translator_slave_araddr),                                          //          .araddr
		.s0_arlen    (axi_translator_slave_arlen),                                           //          .arlen
		.s0_arsize   (axi_translator_slave_arsize),                                          //          .arsize
		.s0_arburst  (axi_translator_slave_arburst),                                         //          .arburst
		.s0_arlock   (axi_translator_slave_arlock),                                          //          .arlock
		.s0_arcache  (axi_translator_slave_arcache),                                         //          .arcache
		.s0_arprot   (axi_translator_slave_arprot),                                          //          .arprot
		.s0_arvalid  (axi_translator_slave_arvalid),                                         //          .arvalid
		.s0_arready  (axi_translator_slave_arready),                                         //          .arready
		.s0_rid      (axi_translator_slave_rid),                                             //          .rid
		.s0_rdata    (axi_translator_slave_rdata),                                           //          .rdata
		.s0_rresp    (axi_translator_slave_rresp),                                           //          .rresp
		.s0_rlast    (axi_translator_slave_rlast),                                           //          .rlast
		.s0_rvalid   (axi_translator_slave_rvalid),                                          //          .rvalid
		.s0_rready   (axi_translator_slave_rready),                                          //          .rready
		.m0_awid     (axi_translator_m0_awid),                                               //        m0.awid
		.m0_awaddr   (axi_translator_m0_awaddr),                                             //          .awaddr
		.m0_awlen    (axi_translator_m0_awlen),                                              //          .awlen
		.m0_awsize   (axi_translator_m0_awsize),                                             //          .awsize
		.m0_awburst  (axi_translator_m0_awburst),                                            //          .awburst
		.m0_awlock   (axi_translator_m0_awlock),                                             //          .awlock
		.m0_awcache  (axi_translator_m0_awcache),                                            //          .awcache
		.m0_awprot   (axi_translator_m0_awprot),                                             //          .awprot
		.m0_awqos    (axi_translator_m0_awqos),                                              //          .awqos
		.m0_awregion (axi_translator_m0_awregion),                                           //          .awregion
		.m0_awvalid  (axi_translator_m0_awvalid),                                            //          .awvalid
		.m0_awready  (axi_translator_m0_awready),                                            //          .awready
		.m0_wdata    (axi_translator_m0_wdata),                                              //          .wdata
		.m0_wstrb    (axi_translator_m0_wstrb),                                              //          .wstrb
		.m0_wlast    (axi_translator_m0_wlast),                                              //          .wlast
		.m0_wvalid   (axi_translator_m0_wvalid),                                             //          .wvalid
		.m0_wready   (axi_translator_m0_wready),                                             //          .wready
		.m0_bid      (axi_translator_m0_bid),                                                //          .bid
		.m0_bresp    (axi_translator_m0_bresp),                                              //          .bresp
		.m0_bvalid   (axi_translator_m0_bvalid),                                             //          .bvalid
		.m0_bready   (axi_translator_m0_bready),                                             //          .bready
		.m0_arid     (axi_translator_m0_arid),                                               //          .arid
		.m0_araddr   (axi_translator_m0_araddr),                                             //          .araddr
		.m0_arlen    (axi_translator_m0_arlen),                                              //          .arlen
		.m0_arsize   (axi_translator_m0_arsize),                                             //          .arsize
		.m0_arburst  (axi_translator_m0_arburst),                                            //          .arburst
		.m0_arlock   (axi_translator_m0_arlock),                                             //          .arlock
		.m0_arcache  (axi_translator_m0_arcache),                                            //          .arcache
		.m0_arprot   (axi_translator_m0_arprot),                                             //          .arprot
		.m0_arqos    (axi_translator_m0_arqos),                                              //          .arqos
		.m0_arregion (axi_translator_m0_arregion),                                           //          .arregion
		.m0_arvalid  (axi_translator_m0_arvalid),                                            //          .arvalid
		.m0_arready  (axi_translator_m0_arready),                                            //          .arready
		.m0_rid      (axi_translator_m0_rid),                                                //          .rid
		.m0_rdata    (axi_translator_m0_rdata),                                              //          .rdata
		.m0_rresp    (axi_translator_m0_rresp),                                              //          .rresp
		.m0_rlast    (axi_translator_m0_rlast),                                              //          .rlast
		.m0_rvalid   (axi_translator_m0_rvalid),                                             //          .rvalid
		.m0_rready   (axi_translator_m0_rready),                                             //          .rready
		.s0_awuser   (64'b0000000000000000000000000000000000000000000000000000000000000000), // (terminated)
		.s0_awqos    (4'b0000),                                                              // (terminated)
		.s0_awregion (4'b0000),                                                              // (terminated)
		.s0_wuser    (64'b0000000000000000000000000000000000000000000000000000000000000000), // (terminated)
		.s0_buser    (),                                                                     // (terminated)
		.s0_aruser   (64'b0000000000000000000000000000000000000000000000000000000000000000), // (terminated)
		.s0_arqos    (4'b0000),                                                              // (terminated)
		.s0_arregion (4'b0000),                                                              // (terminated)
		.s0_ruser    (),                                                                     // (terminated)
		.m0_awuser   (),                                                                     // (terminated)
		.m0_wuser    (),                                                                     // (terminated)
		.m0_buser    (64'b0000000000000000000000000000000000000000000000000000000000000000), // (terminated)
		.m0_aruser   (),                                                                     // (terminated)
		.m0_ruser    (64'b0000000000000000000000000000000000000000000000000000000000000000), // (terminated)
		.s0_wid      (4'b0000),                                                              // (terminated)
		.m0_wid      ()                                                                      // (terminated)
	);

	altera_merlin_axi_translator #(
		.USE_S0_AWID                       (1),
		.USE_S0_AWREGION                   (1),
		.USE_M0_AWREGION                   (1),
		.USE_S0_AWLEN                      (1),
		.USE_S0_AWSIZE                     (1),
		.USE_S0_AWBURST                    (1),
		.USE_S0_AWLOCK                     (1),
		.USE_M0_AWLOCK                     (1),
		.USE_S0_AWCACHE                    (1),
		.USE_M0_AWCACHE                    (1),
		.USE_M0_AWPROT                     (1),
		.USE_S0_AWQOS                      (1),
		.USE_M0_AWQOS                      (1),
		.USE_S0_WSTRB                      (1),
		.USE_M0_WLAST                      (1),
		.USE_S0_BID                        (1),
		.USE_S0_BRESP                      (1),
		.USE_M0_BRESP                      (1),
		.USE_S0_ARID                       (1),
		.USE_S0_ARREGION                   (1),
		.USE_M0_ARREGION                   (1),
		.USE_S0_ARLEN                      (1),
		.USE_S0_ARSIZE                     (1),
		.USE_S0_ARBURST                    (1),
		.USE_S0_ARLOCK                     (1),
		.USE_M0_ARLOCK                     (1),
		.USE_M0_ARCACHE                    (1),
		.USE_M0_ARQOS                      (1),
		.USE_M0_ARPROT                     (1),
		.USE_S0_ARCACHE                    (1),
		.USE_S0_ARQOS                      (1),
		.USE_S0_RID                        (1),
		.USE_S0_RRESP                      (1),
		.USE_M0_RRESP                      (1),
		.USE_S0_RLAST                      (1),
		.M0_ID_WIDTH                       (8),
		.DATA_WIDTH                        (32),
		.S0_ID_WIDTH                       (8),
		.M0_ADDR_WIDTH                     (32),
		.S0_WRITE_ADDR_USER_WIDTH          (1),
		.S0_READ_ADDR_USER_WIDTH           (1),
		.M0_WRITE_ADDR_USER_WIDTH          (1),
		.M0_READ_ADDR_USER_WIDTH           (1),
		.S0_WRITE_DATA_USER_WIDTH          (1),
		.S0_WRITE_RESPONSE_DATA_USER_WIDTH (1),
		.S0_READ_DATA_USER_WIDTH           (1),
		.M0_WRITE_DATA_USER_WIDTH          (1),
		.M0_WRITE_RESPONSE_DATA_USER_WIDTH (1),
		.M0_READ_DATA_USER_WIDTH           (1),
		.S0_ADDR_WIDTH                     (32),
		.USE_S0_AWUSER                     (0),
		.USE_S0_ARUSER                     (0),
		.USE_S0_WUSER                      (0),
		.USE_S0_RUSER                      (0),
		.USE_S0_BUSER                      (0),
		.USE_M0_AWUSER                     (1),
		.USE_M0_ARUSER                     (1),
		.USE_M0_WUSER                      (1),
		.USE_M0_RUSER                      (1),
		.USE_M0_BUSER                      (1),
		.M0_AXI_VERSION                    ("AXI4"),
		.M0_BURST_LENGTH_WIDTH             (8),
		.S0_BURST_LENGTH_WIDTH             (8),
		.M0_LOCK_WIDTH                     (1),
		.S0_LOCK_WIDTH                     (1),
		.S0_AXI_VERSION                    ("AXI4")
	) axi_translator_m0_translator (
		.aclk        (clk_clk),                                  //       clk.clk
		.aresetn     (~rst_controller_reset_out_reset),          // clk_reset.reset_n
		.s0_awid     (axi_translator_m0_awid),                   //        s0.awid
		.s0_awaddr   (axi_translator_m0_awaddr),                 //          .awaddr
		.s0_awlen    (axi_translator_m0_awlen),                  //          .awlen
		.s0_awsize   (axi_translator_m0_awsize),                 //          .awsize
		.s0_awburst  (axi_translator_m0_awburst),                //          .awburst
		.s0_awlock   (axi_translator_m0_awlock),                 //          .awlock
		.s0_awcache  (axi_translator_m0_awcache),                //          .awcache
		.s0_awprot   (axi_translator_m0_awprot),                 //          .awprot
		.s0_awqos    (axi_translator_m0_awqos),                  //          .awqos
		.s0_awregion (axi_translator_m0_awregion),               //          .awregion
		.s0_awvalid  (axi_translator_m0_awvalid),                //          .awvalid
		.s0_awready  (axi_translator_m0_awready),                //          .awready
		.s0_wdata    (axi_translator_m0_wdata),                  //          .wdata
		.s0_wstrb    (axi_translator_m0_wstrb),                  //          .wstrb
		.s0_wlast    (axi_translator_m0_wlast),                  //          .wlast
		.s0_wvalid   (axi_translator_m0_wvalid),                 //          .wvalid
		.s0_wready   (axi_translator_m0_wready),                 //          .wready
		.s0_bid      (axi_translator_m0_bid),                    //          .bid
		.s0_bresp    (axi_translator_m0_bresp),                  //          .bresp
		.s0_bvalid   (axi_translator_m0_bvalid),                 //          .bvalid
		.s0_bready   (axi_translator_m0_bready),                 //          .bready
		.s0_arid     (axi_translator_m0_arid),                   //          .arid
		.s0_araddr   (axi_translator_m0_araddr),                 //          .araddr
		.s0_arlen    (axi_translator_m0_arlen),                  //          .arlen
		.s0_arsize   (axi_translator_m0_arsize),                 //          .arsize
		.s0_arburst  (axi_translator_m0_arburst),                //          .arburst
		.s0_arlock   (axi_translator_m0_arlock),                 //          .arlock
		.s0_arcache  (axi_translator_m0_arcache),                //          .arcache
		.s0_arprot   (axi_translator_m0_arprot),                 //          .arprot
		.s0_arqos    (axi_translator_m0_arqos),                  //          .arqos
		.s0_arregion (axi_translator_m0_arregion),               //          .arregion
		.s0_arvalid  (axi_translator_m0_arvalid),                //          .arvalid
		.s0_arready  (axi_translator_m0_arready),                //          .arready
		.s0_rid      (axi_translator_m0_rid),                    //          .rid
		.s0_rdata    (axi_translator_m0_rdata),                  //          .rdata
		.s0_rresp    (axi_translator_m0_rresp),                  //          .rresp
		.s0_rlast    (axi_translator_m0_rlast),                  //          .rlast
		.s0_rvalid   (axi_translator_m0_rvalid),                 //          .rvalid
		.s0_rready   (axi_translator_m0_rready),                 //          .rready
		.m0_awid     (axi_translator_m0_translator_m0_awid),     //        m0.awid
		.m0_awaddr   (axi_translator_m0_translator_m0_awaddr),   //          .awaddr
		.m0_awlen    (axi_translator_m0_translator_m0_awlen),    //          .awlen
		.m0_awsize   (axi_translator_m0_translator_m0_awsize),   //          .awsize
		.m0_awburst  (axi_translator_m0_translator_m0_awburst),  //          .awburst
		.m0_awlock   (axi_translator_m0_translator_m0_awlock),   //          .awlock
		.m0_awcache  (axi_translator_m0_translator_m0_awcache),  //          .awcache
		.m0_awprot   (axi_translator_m0_translator_m0_awprot),   //          .awprot
		.m0_awuser   (axi_translator_m0_translator_m0_awuser),   //          .awuser
		.m0_awqos    (axi_translator_m0_translator_m0_awqos),    //          .awqos
		.m0_awregion (axi_translator_m0_translator_m0_awregion), //          .awregion
		.m0_awvalid  (axi_translator_m0_translator_m0_awvalid),  //          .awvalid
		.m0_awready  (axi_translator_m0_translator_m0_awready),  //          .awready
		.m0_wdata    (axi_translator_m0_translator_m0_wdata),    //          .wdata
		.m0_wstrb    (axi_translator_m0_translator_m0_wstrb),    //          .wstrb
		.m0_wlast    (axi_translator_m0_translator_m0_wlast),    //          .wlast
		.m0_wvalid   (axi_translator_m0_translator_m0_wvalid),   //          .wvalid
		.m0_wuser    (axi_translator_m0_translator_m0_wuser),    //          .wuser
		.m0_wready   (axi_translator_m0_translator_m0_wready),   //          .wready
		.m0_bid      (axi_translator_m0_translator_m0_bid),      //          .bid
		.m0_bresp    (axi_translator_m0_translator_m0_bresp),    //          .bresp
		.m0_buser    (axi_translator_m0_translator_m0_buser),    //          .buser
		.m0_bvalid   (axi_translator_m0_translator_m0_bvalid),   //          .bvalid
		.m0_bready   (axi_translator_m0_translator_m0_bready),   //          .bready
		.m0_arid     (axi_translator_m0_translator_m0_arid),     //          .arid
		.m0_araddr   (axi_translator_m0_translator_m0_araddr),   //          .araddr
		.m0_arlen    (axi_translator_m0_translator_m0_arlen),    //          .arlen
		.m0_arsize   (axi_translator_m0_translator_m0_arsize),   //          .arsize
		.m0_arburst  (axi_translator_m0_translator_m0_arburst),  //          .arburst
		.m0_arlock   (axi_translator_m0_translator_m0_arlock),   //          .arlock
		.m0_arcache  (axi_translator_m0_translator_m0_arcache),  //          .arcache
		.m0_arprot   (axi_translator_m0_translator_m0_arprot),   //          .arprot
		.m0_aruser   (axi_translator_m0_translator_m0_aruser),   //          .aruser
		.m0_arqos    (axi_translator_m0_translator_m0_arqos),    //          .arqos
		.m0_arregion (axi_translator_m0_translator_m0_arregion), //          .arregion
		.m0_arvalid  (axi_translator_m0_translator_m0_arvalid),  //          .arvalid
		.m0_arready  (axi_translator_m0_translator_m0_arready),  //          .arready
		.m0_rid      (axi_translator_m0_translator_m0_rid),      //          .rid
		.m0_rdata    (axi_translator_m0_translator_m0_rdata),    //          .rdata
		.m0_rresp    (axi_translator_m0_translator_m0_rresp),    //          .rresp
		.m0_rlast    (axi_translator_m0_translator_m0_rlast),    //          .rlast
		.m0_rvalid   (axi_translator_m0_translator_m0_rvalid),   //          .rvalid
		.m0_rready   (axi_translator_m0_translator_m0_rready),   //          .rready
		.m0_ruser    (axi_translator_m0_translator_m0_ruser),    //          .ruser
		.s0_awuser   (1'b0),                                     // (terminated)
		.s0_wuser    (1'b0),                                     // (terminated)
		.s0_buser    (),                                         // (terminated)
		.s0_aruser   (1'b0),                                     // (terminated)
		.s0_ruser    (),                                         // (terminated)
		.s0_wid      (8'b00000000),                              // (terminated)
		.m0_wid      ()                                          // (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (24),
		.AV_DATA_W                      (128),
		.UAV_DATA_W                     (128),
		.AV_BURSTCOUNT_W                (6),
		.AV_BYTEENABLE_W                (16),
		.UAV_BYTEENABLE_W               (16),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (10),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (16),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mem_if_ddr3_emif_0_avl_translator (
		.clk                      (mem_if_ddr3_emif_0_afi_clk_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                //                    reset.reset
		.uav_address              (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_beginbursttransfer    (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_beginbursttransfer),          //                         .beginbursttransfer
		.av_burstcount            (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (~mem_if_ddr3_emif_0_avl_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_chipselect            (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_axi_master_ni #(
		.ID_WIDTH                  (8),
		.ADDR_WIDTH                (32),
		.RDATA_WIDTH               (32),
		.WDATA_WIDTH               (32),
		.ADDR_USER_WIDTH           (1),
		.DATA_USER_WIDTH           (1),
		.AXI_BURST_LENGTH_WIDTH    (8),
		.AXI_LOCK_WIDTH            (1),
		.AXI_VERSION               ("AXI4"),
		.WRITE_ISSUING_CAPABILITY  (16),
		.READ_ISSUING_CAPABILITY   (16),
		.PKT_BEGIN_BURST           (101),
		.PKT_CACHE_H               (122),
		.PKT_CACHE_L               (119),
		.PKT_ADDR_SIDEBAND_H       (99),
		.PKT_ADDR_SIDEBAND_L       (99),
		.PKT_PROTECTION_H          (118),
		.PKT_PROTECTION_L          (116),
		.PKT_BURST_SIZE_H          (96),
		.PKT_BURST_SIZE_L          (94),
		.PKT_BURST_TYPE_H          (98),
		.PKT_BURST_TYPE_L          (97),
		.PKT_RESPONSE_STATUS_L     (123),
		.PKT_RESPONSE_STATUS_H     (124),
		.PKT_BURSTWRAP_H           (93),
		.PKT_BURSTWRAP_L           (87),
		.PKT_BYTE_CNT_H            (86),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (106),
		.PKT_SRC_ID_L              (106),
		.PKT_DEST_ID_H             (107),
		.PKT_DEST_ID_L             (107),
		.PKT_THREAD_ID_H           (115),
		.PKT_THREAD_ID_L           (108),
		.PKT_QOS_L                 (102),
		.PKT_QOS_H                 (105),
		.PKT_DATA_SIDEBAND_H       (100),
		.PKT_DATA_SIDEBAND_L       (100),
		.ST_DATA_W                 (125),
		.ST_CHANNEL_W              (2),
		.ID                        (0)
	) axi_translator_m0_translator_m0_agent (
		.aclk                   (clk_clk),                                                      //              clk.clk
		.aresetn                (~rst_controller_reset_out_reset),                              //        clk_reset.reset_n
		.write_cp_valid         (axi_translator_m0_translator_m0_agent_write_cp_valid),         //         write_cp.valid
		.write_cp_data          (axi_translator_m0_translator_m0_agent_write_cp_data),          //                 .data
		.write_cp_startofpacket (axi_translator_m0_translator_m0_agent_write_cp_startofpacket), //                 .startofpacket
		.write_cp_endofpacket   (axi_translator_m0_translator_m0_agent_write_cp_endofpacket),   //                 .endofpacket
		.write_cp_ready         (axi_translator_m0_translator_m0_agent_write_cp_ready),         //                 .ready
		.write_rp_valid         (crosser_002_out_valid),                                        //         write_rp.valid
		.write_rp_data          (crosser_002_out_data),                                         //                 .data
		.write_rp_channel       (crosser_002_out_channel),                                      //                 .channel
		.write_rp_startofpacket (crosser_002_out_startofpacket),                                //                 .startofpacket
		.write_rp_endofpacket   (crosser_002_out_endofpacket),                                  //                 .endofpacket
		.write_rp_ready         (crosser_002_out_ready),                                        //                 .ready
		.read_cp_valid          (axi_translator_m0_translator_m0_agent_read_cp_valid),          //          read_cp.valid
		.read_cp_data           (axi_translator_m0_translator_m0_agent_read_cp_data),           //                 .data
		.read_cp_startofpacket  (axi_translator_m0_translator_m0_agent_read_cp_startofpacket),  //                 .startofpacket
		.read_cp_endofpacket    (axi_translator_m0_translator_m0_agent_read_cp_endofpacket),    //                 .endofpacket
		.read_cp_ready          (axi_translator_m0_translator_m0_agent_read_cp_ready),          //                 .ready
		.read_rp_valid          (crosser_003_out_valid),                                        //          read_rp.valid
		.read_rp_data           (crosser_003_out_data),                                         //                 .data
		.read_rp_channel        (crosser_003_out_channel),                                      //                 .channel
		.read_rp_startofpacket  (crosser_003_out_startofpacket),                                //                 .startofpacket
		.read_rp_endofpacket    (crosser_003_out_endofpacket),                                  //                 .endofpacket
		.read_rp_ready          (crosser_003_out_ready),                                        //                 .ready
		.awid                   (axi_translator_m0_translator_m0_awid),                         // altera_axi_slave.awid
		.awaddr                 (axi_translator_m0_translator_m0_awaddr),                       //                 .awaddr
		.awlen                  (axi_translator_m0_translator_m0_awlen),                        //                 .awlen
		.awsize                 (axi_translator_m0_translator_m0_awsize),                       //                 .awsize
		.awburst                (axi_translator_m0_translator_m0_awburst),                      //                 .awburst
		.awlock                 (axi_translator_m0_translator_m0_awlock),                       //                 .awlock
		.awcache                (axi_translator_m0_translator_m0_awcache),                      //                 .awcache
		.awprot                 (axi_translator_m0_translator_m0_awprot),                       //                 .awprot
		.awuser                 (axi_translator_m0_translator_m0_awuser),                       //                 .awuser
		.awqos                  (axi_translator_m0_translator_m0_awqos),                        //                 .awqos
		.awregion               (axi_translator_m0_translator_m0_awregion),                     //                 .awregion
		.awvalid                (axi_translator_m0_translator_m0_awvalid),                      //                 .awvalid
		.awready                (axi_translator_m0_translator_m0_awready),                      //                 .awready
		.wdata                  (axi_translator_m0_translator_m0_wdata),                        //                 .wdata
		.wstrb                  (axi_translator_m0_translator_m0_wstrb),                        //                 .wstrb
		.wlast                  (axi_translator_m0_translator_m0_wlast),                        //                 .wlast
		.wvalid                 (axi_translator_m0_translator_m0_wvalid),                       //                 .wvalid
		.wuser                  (axi_translator_m0_translator_m0_wuser),                        //                 .wuser
		.wready                 (axi_translator_m0_translator_m0_wready),                       //                 .wready
		.bid                    (axi_translator_m0_translator_m0_bid),                          //                 .bid
		.bresp                  (axi_translator_m0_translator_m0_bresp),                        //                 .bresp
		.buser                  (axi_translator_m0_translator_m0_buser),                        //                 .buser
		.bvalid                 (axi_translator_m0_translator_m0_bvalid),                       //                 .bvalid
		.bready                 (axi_translator_m0_translator_m0_bready),                       //                 .bready
		.arid                   (axi_translator_m0_translator_m0_arid),                         //                 .arid
		.araddr                 (axi_translator_m0_translator_m0_araddr),                       //                 .araddr
		.arlen                  (axi_translator_m0_translator_m0_arlen),                        //                 .arlen
		.arsize                 (axi_translator_m0_translator_m0_arsize),                       //                 .arsize
		.arburst                (axi_translator_m0_translator_m0_arburst),                      //                 .arburst
		.arlock                 (axi_translator_m0_translator_m0_arlock),                       //                 .arlock
		.arcache                (axi_translator_m0_translator_m0_arcache),                      //                 .arcache
		.arprot                 (axi_translator_m0_translator_m0_arprot),                       //                 .arprot
		.aruser                 (axi_translator_m0_translator_m0_aruser),                       //                 .aruser
		.arqos                  (axi_translator_m0_translator_m0_arqos),                        //                 .arqos
		.arregion               (axi_translator_m0_translator_m0_arregion),                     //                 .arregion
		.arvalid                (axi_translator_m0_translator_m0_arvalid),                      //                 .arvalid
		.arready                (axi_translator_m0_translator_m0_arready),                      //                 .arready
		.rid                    (axi_translator_m0_translator_m0_rid),                          //                 .rid
		.rdata                  (axi_translator_m0_translator_m0_rdata),                        //                 .rdata
		.rresp                  (axi_translator_m0_translator_m0_rresp),                        //                 .rresp
		.rlast                  (axi_translator_m0_translator_m0_rlast),                        //                 .rlast
		.rvalid                 (axi_translator_m0_translator_m0_rvalid),                       //                 .rvalid
		.rready                 (axi_translator_m0_translator_m0_rready),                       //                 .rready
		.ruser                  (axi_translator_m0_translator_m0_ruser),                        //                 .ruser
		.wid                    (8'b00000000)                                                   //      (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (127),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (209),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (143),
		.PKT_BYTEEN_L              (128),
		.PKT_ADDR_H                (175),
		.PKT_ADDR_L                (144),
		.PKT_TRANS_COMPRESSED_READ (176),
		.PKT_TRANS_POSTED          (177),
		.PKT_TRANS_WRITE           (178),
		.PKT_TRANS_READ            (179),
		.PKT_TRANS_LOCK            (180),
		.PKT_SRC_ID_H              (214),
		.PKT_SRC_ID_L              (214),
		.PKT_DEST_ID_H             (215),
		.PKT_DEST_ID_L             (215),
		.PKT_BURSTWRAP_H           (201),
		.PKT_BURSTWRAP_L           (195),
		.PKT_BYTE_CNT_H            (194),
		.PKT_BYTE_CNT_L            (182),
		.PKT_PROTECTION_H          (226),
		.PKT_PROTECTION_L          (224),
		.PKT_RESPONSE_STATUS_H     (232),
		.PKT_RESPONSE_STATUS_L     (231),
		.PKT_BURST_SIZE_H          (204),
		.PKT_BURST_SIZE_L          (202),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (233),
		.AVS_BURSTCOUNT_W          (10),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent (
		.clk                     (mem_if_ddr3_emif_0_afi_clk_clk),                                                              //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                                 //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                                 //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                  //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                           //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                               //                .channel
		.rf_sink_ready           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (234),
		.FIFO_DEPTH          (33),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (mem_if_ddr3_emif_0_afi_clk_clk),                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (130),
		.FIFO_DEPTH          (2048),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (mem_if_ddr3_emif_0_afi_clk_clk),                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_startofpacket  (1'b0),                                                                                  // (terminated)
		.in_endofpacket    (1'b0),                                                                                  // (terminated)
		.out_startofpacket (),                                                                                      // (terminated)
		.out_endofpacket   (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	fpga_sdram_controller_addr_router addr_router (
		.sink_ready         (axi_translator_m0_translator_m0_agent_write_cp_ready),         //      sink.ready
		.sink_valid         (axi_translator_m0_translator_m0_agent_write_cp_valid),         //          .valid
		.sink_data          (axi_translator_m0_translator_m0_agent_write_cp_data),          //          .data
		.sink_startofpacket (axi_translator_m0_translator_m0_agent_write_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (axi_translator_m0_translator_m0_agent_write_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                               // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                        //       src.ready
		.src_valid          (addr_router_src_valid),                                        //          .valid
		.src_data           (addr_router_src_data),                                         //          .data
		.src_channel        (addr_router_src_channel),                                      //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                   //          .endofpacket
	);

	fpga_sdram_controller_addr_router addr_router_001 (
		.sink_ready         (axi_translator_m0_translator_m0_agent_read_cp_ready),         //      sink.ready
		.sink_valid         (axi_translator_m0_translator_m0_agent_read_cp_valid),         //          .valid
		.sink_data          (axi_translator_m0_translator_m0_agent_read_cp_data),          //          .data
		.sink_startofpacket (axi_translator_m0_translator_m0_agent_read_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (axi_translator_m0_translator_m0_agent_read_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                              // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                   //       src.ready
		.src_valid          (addr_router_001_src_valid),                                   //          .valid
		.src_data           (addr_router_001_src_data),                                    //          .data
		.src_channel        (addr_router_001_src_channel),                                 //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                           //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                              //          .endofpacket
	);

	fpga_sdram_controller_id_router id_router (
		.sink_ready         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mem_if_ddr3_emif_0_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (mem_if_ddr3_emif_0_afi_clk_clk),                                                    //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                               //       src.ready
		.src_valid          (id_router_src_valid),                                                               //          .valid
		.src_data           (id_router_src_data),                                                                //          .data
		.src_channel        (id_router_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                          //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (175),
		.PKT_ADDR_L                (144),
		.PKT_BEGIN_BURST           (209),
		.PKT_BYTE_CNT_H            (194),
		.PKT_BYTE_CNT_L            (182),
		.PKT_BYTEEN_H              (143),
		.PKT_BYTEEN_L              (128),
		.PKT_BURST_SIZE_H          (204),
		.PKT_BURST_SIZE_L          (202),
		.PKT_BURST_TYPE_H          (206),
		.PKT_BURST_TYPE_L          (205),
		.PKT_BURSTWRAP_H           (201),
		.PKT_BURSTWRAP_L           (195),
		.PKT_TRANS_COMPRESSED_READ (176),
		.PKT_TRANS_WRITE           (178),
		.PKT_TRANS_READ            (179),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (1),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (233),
		.ST_CHANNEL_W              (2),
		.OUT_BYTE_CNT_H            (191),
		.OUT_BURSTWRAP_H           (201),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (0),
		.BURSTWRAP_CONST_VALUE     (0)
	) burst_adapter (
		.clk                   (mem_if_ddr3_emif_0_afi_clk_clk),         //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),     // cr0_reset.reset
		.sink0_valid           (width_adapter_cmd_source_valid),         //     sink0.valid
		.sink0_data            (width_adapter_cmd_source_data),          //          .data
		.sink0_channel         (width_adapter_cmd_source_channel),       //          .channel
		.sink0_startofpacket   (width_adapter_cmd_source_startofpacket), //          .startofpacket
		.sink0_endofpacket     (width_adapter_cmd_source_endofpacket),   //          .endofpacket
		.sink0_ready           (width_adapter_cmd_source_ready),         //          .ready
		.source0_valid         (burst_adapter_source0_valid),            //   source0.valid
		.source0_data          (burst_adapter_source0_data),             //          .data
		.source0_channel       (burst_adapter_source0_channel),          //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket),    //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),      //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)             //          .ready
	);

	altera_merlin_combined_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (86),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (93),
		.IN_PKT_BURSTWRAP_L            (87),
		.IN_PKT_BURST_SIZE_H           (96),
		.IN_PKT_BURST_SIZE_L           (94),
		.IN_PKT_RESPONSE_STATUS_H      (124),
		.IN_PKT_RESPONSE_STATUS_L      (123),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (98),
		.IN_PKT_BURST_TYPE_L           (97),
		.IN_PKT_TRANS_POSTED           (69),
		.IN_ST_DATA_W                  (125),
		.OUT_PKT_ADDR_H                (175),
		.OUT_PKT_ADDR_L                (144),
		.OUT_PKT_DATA_H                (127),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (143),
		.OUT_PKT_BYTEEN_L              (128),
		.OUT_PKT_BYTE_CNT_H            (194),
		.OUT_PKT_BYTE_CNT_L            (182),
		.OUT_PKT_TRANS_COMPRESSED_READ (176),
		.OUT_PKT_TRANS_EXCLUSIVE       (181),
		.OUT_PKT_RESPONSE_STATUS_H     (232),
		.OUT_PKT_RESPONSE_STATUS_L     (231),
		.OUT_PKT_BURST_SIZE_H          (204),
		.OUT_PKT_BURST_SIZE_L          (202),
		.OUT_PKT_BURST_TYPE_H          (206),
		.OUT_PKT_BURST_TYPE_L          (205),
		.OUT_ST_DATA_W                 (233),
		.ST_CHANNEL_W                  (2),
		.MAX_OUTSTANDING_RESPONSES     (40)
	) width_adapter (
		.clk                   (mem_if_ddr3_emif_0_afi_clk_clk),         //      clock.clk
		.reset                 (rst_controller_001_reset_out_reset),     //      reset.reset
		.cmd_in_valid          (cmd_xbar_mux_src_valid),                 //   cmd_sink.valid
		.cmd_in_channel        (cmd_xbar_mux_src_channel),               //           .channel
		.cmd_in_data           (cmd_xbar_mux_src_data),                  //           .data
		.cmd_in_startofpacket  (cmd_xbar_mux_src_startofpacket),         //           .startofpacket
		.cmd_in_endofpacket    (cmd_xbar_mux_src_endofpacket),           //           .endofpacket
		.cmd_in_ready          (cmd_xbar_mux_src_ready),                 //           .ready
		.cmd_out_ready         (width_adapter_cmd_source_ready),         // cmd_source.ready
		.cmd_out_valid         (width_adapter_cmd_source_valid),         //           .valid
		.cmd_out_channel       (width_adapter_cmd_source_channel),       //           .channel
		.cmd_out_data          (width_adapter_cmd_source_data),          //           .data
		.cmd_out_startofpacket (width_adapter_cmd_source_startofpacket), //           .startofpacket
		.cmd_out_endofpacket   (width_adapter_cmd_source_endofpacket),   //           .endofpacket
		.rsp_in_ready          (id_router_src_ready),                    //   rsp_sink.ready
		.rsp_in_valid          (id_router_src_valid),                    //           .valid
		.rsp_in_channel        (id_router_src_channel),                  //           .channel
		.rsp_in_data           (id_router_src_data),                     //           .data
		.rsp_in_startofpacket  (id_router_src_startofpacket),            //           .startofpacket
		.rsp_in_endofpacket    (id_router_src_endofpacket),              //           .endofpacket
		.rsp_out_ready         (width_adapter_rsp_source_ready),         // rsp_source.ready
		.rsp_out_valid         (width_adapter_rsp_source_valid),         //           .valid
		.rsp_out_channel       (width_adapter_rsp_source_channel),       //           .channel
		.rsp_out_data          (width_adapter_rsp_source_data),          //           .data
		.rsp_out_startofpacket (width_adapter_rsp_source_startofpacket), //           .startofpacket
		.rsp_out_endofpacket   (width_adapter_rsp_source_endofpacket)    //           .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~mem_if_ddr3_emif_0_afi_reset_reset), // reset_in0.reset
		.clk        (mem_if_ddr3_emif_0_afi_clk_clk),      //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_req  (),                                    // (terminated)
		.reset_in1  (1'b0),                                // (terminated)
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	fpga_sdram_controller_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	fpga_sdram_controller_cmd_xbar_demux cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	fpga_sdram_controller_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (mem_if_ddr3_emif_0_afi_clk_clk),     //       clk.clk
		.reset               (rst_controller_001_reset_out_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),       //          .endofpacket
		.sink0_ready         (crosser_out_ready),                  //     sink0.ready
		.sink0_valid         (crosser_out_valid),                  //          .valid
		.sink0_channel       (crosser_out_channel),                //          .channel
		.sink0_data          (crosser_out_data),                   //          .data
		.sink0_startofpacket (crosser_out_startofpacket),          //          .startofpacket
		.sink0_endofpacket   (crosser_out_endofpacket),            //          .endofpacket
		.sink1_ready         (crosser_001_out_ready),              //     sink1.ready
		.sink1_valid         (crosser_001_out_valid),              //          .valid
		.sink1_channel       (crosser_001_out_channel),            //          .channel
		.sink1_data          (crosser_001_out_data),               //          .data
		.sink1_startofpacket (crosser_001_out_startofpacket),      //          .startofpacket
		.sink1_endofpacket   (crosser_001_out_endofpacket)         //          .endofpacket
	);

	fpga_sdram_controller_rsp_xbar_demux rsp_xbar_demux (
		.clk                (mem_if_ddr3_emif_0_afi_clk_clk),         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.sink_ready         (width_adapter_rsp_source_ready),         //      sink.ready
		.sink_channel       (width_adapter_rsp_source_channel),       //          .channel
		.sink_data          (width_adapter_rsp_source_data),          //          .data
		.sink_startofpacket (width_adapter_rsp_source_startofpacket), //          .startofpacket
		.sink_endofpacket   (width_adapter_rsp_source_endofpacket),   //          .endofpacket
		.sink_valid         (width_adapter_rsp_source_valid),         //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),              //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),              //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),               //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),            //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),      //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),        //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),              //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),              //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),               //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),            //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),      //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)         //          .endofpacket
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (125),
		.BITS_PER_SYMBOL     (125),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (2),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (clk_clk),                            //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),     //  in_clk_reset.reset
		.out_clk           (mem_if_ddr3_emif_0_afi_clk_clk),     //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset), // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src0_ready),          //            in.ready
		.in_valid          (cmd_xbar_demux_src0_valid),          //              .valid
		.in_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //              .endofpacket
		.in_channel        (cmd_xbar_demux_src0_channel),        //              .channel
		.in_data           (cmd_xbar_demux_src0_data),           //              .data
		.out_ready         (crosser_out_ready),                  //           out.ready
		.out_valid         (crosser_out_valid),                  //              .valid
		.out_startofpacket (crosser_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_out_channel),                //              .channel
		.out_data          (crosser_out_data),                   //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (125),
		.BITS_PER_SYMBOL     (125),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (2),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (mem_if_ddr3_emif_0_afi_clk_clk),        //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (125),
		.BITS_PER_SYMBOL     (125),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (2),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (mem_if_ddr3_emif_0_afi_clk_clk),     //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset), //  in_clk_reset.reset
		.out_clk           (clk_clk),                            //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_src0_ready),          //            in.ready
		.in_valid          (rsp_xbar_demux_src0_valid),          //              .valid
		.in_startofpacket  (rsp_xbar_demux_src0_startofpacket),  //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_src0_endofpacket),    //              .endofpacket
		.in_channel        (rsp_xbar_demux_src0_channel),        //              .channel
		.in_data           (rsp_xbar_demux_src0_data),           //              .data
		.out_ready         (crosser_002_out_ready),              //           out.ready
		.out_valid         (crosser_002_out_valid),              //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),      //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),        //              .endofpacket
		.out_channel       (crosser_002_out_channel),            //              .channel
		.out_data          (crosser_002_out_data),               //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (125),
		.BITS_PER_SYMBOL     (125),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (2),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (mem_if_ddr3_emif_0_afi_clk_clk),     //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset), //  in_clk_reset.reset
		.out_clk           (clk_clk),                            //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_src1_ready),          //            in.ready
		.in_valid          (rsp_xbar_demux_src1_valid),          //              .valid
		.in_startofpacket  (rsp_xbar_demux_src1_startofpacket),  //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_src1_endofpacket),    //              .endofpacket
		.in_channel        (rsp_xbar_demux_src1_channel),        //              .channel
		.in_data           (rsp_xbar_demux_src1_data),           //              .data
		.out_ready         (crosser_003_out_ready),              //           out.ready
		.out_valid         (crosser_003_out_valid),              //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),      //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),        //              .endofpacket
		.out_channel       (crosser_003_out_channel),            //              .channel
		.out_data          (crosser_003_out_data),               //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

endmodule
