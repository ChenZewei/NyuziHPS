// HPS.v

// Generated using ACDS version 13.0sp1 232 at 2015.08.07.21:19:15

`timescale 1 ps / 1 ps
module HPS (
		input  wire        clk_clk,            //        clk.clk
		input  wire        reset_reset_n,      //      reset.reset_n
		output wire [12:0] memory_mem_a,       //     memory.mem_a
		output wire [2:0]  memory_mem_ba,      //           .mem_ba
		output wire        memory_mem_ck,      //           .mem_ck
		output wire        memory_mem_ck_n,    //           .mem_ck_n
		output wire        memory_mem_cke,     //           .mem_cke
		output wire        memory_mem_cs_n,    //           .mem_cs_n
		output wire        memory_mem_ras_n,   //           .mem_ras_n
		output wire        memory_mem_cas_n,   //           .mem_cas_n
		output wire        memory_mem_we_n,    //           .mem_we_n
		output wire        memory_mem_reset_n, //           .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,      //           .mem_dq
		inout  wire        memory_mem_dqs,     //           .mem_dqs
		inout  wire        memory_mem_dqs_n,   //           .mem_dqs_n
		output wire        memory_mem_odt,     //           .mem_odt
		output wire        memory_mem_dm,      //           .mem_dm
		input  wire        memory_oct_rzqin,   //           .oct_rzqin
		output wire [11:0] axi_master_awid,    // axi_master.awid
		output wire [29:0] axi_master_awaddr,  //           .awaddr
		output wire [3:0]  axi_master_awlen,   //           .awlen
		output wire [2:0]  axi_master_awsize,  //           .awsize
		output wire [1:0]  axi_master_awburst, //           .awburst
		output wire [1:0]  axi_master_awlock,  //           .awlock
		output wire [3:0]  axi_master_awcache, //           .awcache
		output wire [2:0]  axi_master_awprot,  //           .awprot
		output wire        axi_master_awvalid, //           .awvalid
		input  wire        axi_master_awready, //           .awready
		output wire [11:0] axi_master_wid,     //           .wid
		output wire [63:0] axi_master_wdata,   //           .wdata
		output wire [7:0]  axi_master_wstrb,   //           .wstrb
		output wire        axi_master_wlast,   //           .wlast
		output wire        axi_master_wvalid,  //           .wvalid
		input  wire        axi_master_wready,  //           .wready
		input  wire [11:0] axi_master_bid,     //           .bid
		input  wire [1:0]  axi_master_bresp,   //           .bresp
		input  wire        axi_master_bvalid,  //           .bvalid
		output wire        axi_master_bready,  //           .bready
		output wire [11:0] axi_master_arid,    //           .arid
		output wire [29:0] axi_master_araddr,  //           .araddr
		output wire [3:0]  axi_master_arlen,   //           .arlen
		output wire [2:0]  axi_master_arsize,  //           .arsize
		output wire [1:0]  axi_master_arburst, //           .arburst
		output wire [1:0]  axi_master_arlock,  //           .arlock
		output wire [3:0]  axi_master_arcache, //           .arcache
		output wire [2:0]  axi_master_arprot,  //           .arprot
		output wire        axi_master_arvalid, //           .arvalid
		input  wire        axi_master_arready, //           .arready
		input  wire [11:0] axi_master_rid,     //           .rid
		input  wire [63:0] axi_master_rdata,   //           .rdata
		input  wire [1:0]  axi_master_rresp,   //           .rresp
		input  wire        axi_master_rlast,   //           .rlast
		input  wire        axi_master_rvalid,  //           .rvalid
		output wire        axi_master_rready   //           .rready
	);

	HPS_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (2)
	) hps_0 (
		.mem_a       (memory_mem_a),       //         memory.mem_a
		.mem_ba      (memory_mem_ba),      //               .mem_ba
		.mem_ck      (memory_mem_ck),      //               .mem_ck
		.mem_ck_n    (memory_mem_ck_n),    //               .mem_ck_n
		.mem_cke     (memory_mem_cke),     //               .mem_cke
		.mem_cs_n    (memory_mem_cs_n),    //               .mem_cs_n
		.mem_ras_n   (memory_mem_ras_n),   //               .mem_ras_n
		.mem_cas_n   (memory_mem_cas_n),   //               .mem_cas_n
		.mem_we_n    (memory_mem_we_n),    //               .mem_we_n
		.mem_reset_n (memory_mem_reset_n), //               .mem_reset_n
		.mem_dq      (memory_mem_dq),      //               .mem_dq
		.mem_dqs     (memory_mem_dqs),     //               .mem_dqs
		.mem_dqs_n   (memory_mem_dqs_n),   //               .mem_dqs_n
		.mem_odt     (memory_mem_odt),     //               .mem_odt
		.mem_dm      (memory_mem_dm),      //               .mem_dm
		.oct_rzqin   (memory_oct_rzqin),   //               .oct_rzqin
		.h2f_rst_n   (),                   //      h2f_reset.reset_n
		.h2f_axi_clk (clk_clk),            //  h2f_axi_clock.clk
		.h2f_AWID    (axi_master_awid),    // h2f_axi_master.awid
		.h2f_AWADDR  (axi_master_awaddr),  //               .awaddr
		.h2f_AWLEN   (axi_master_awlen),   //               .awlen
		.h2f_AWSIZE  (axi_master_awsize),  //               .awsize
		.h2f_AWBURST (axi_master_awburst), //               .awburst
		.h2f_AWLOCK  (axi_master_awlock),  //               .awlock
		.h2f_AWCACHE (axi_master_awcache), //               .awcache
		.h2f_AWPROT  (axi_master_awprot),  //               .awprot
		.h2f_AWVALID (axi_master_awvalid), //               .awvalid
		.h2f_AWREADY (axi_master_awready), //               .awready
		.h2f_WID     (axi_master_wid),     //               .wid
		.h2f_WDATA   (axi_master_wdata),   //               .wdata
		.h2f_WSTRB   (axi_master_wstrb),   //               .wstrb
		.h2f_WLAST   (axi_master_wlast),   //               .wlast
		.h2f_WVALID  (axi_master_wvalid),  //               .wvalid
		.h2f_WREADY  (axi_master_wready),  //               .wready
		.h2f_BID     (axi_master_bid),     //               .bid
		.h2f_BRESP   (axi_master_bresp),   //               .bresp
		.h2f_BVALID  (axi_master_bvalid),  //               .bvalid
		.h2f_BREADY  (axi_master_bready),  //               .bready
		.h2f_ARID    (axi_master_arid),    //               .arid
		.h2f_ARADDR  (axi_master_araddr),  //               .araddr
		.h2f_ARLEN   (axi_master_arlen),   //               .arlen
		.h2f_ARSIZE  (axi_master_arsize),  //               .arsize
		.h2f_ARBURST (axi_master_arburst), //               .arburst
		.h2f_ARLOCK  (axi_master_arlock),  //               .arlock
		.h2f_ARCACHE (axi_master_arcache), //               .arcache
		.h2f_ARPROT  (axi_master_arprot),  //               .arprot
		.h2f_ARVALID (axi_master_arvalid), //               .arvalid
		.h2f_ARREADY (axi_master_arready), //               .arready
		.h2f_RID     (axi_master_rid),     //               .rid
		.h2f_RDATA   (axi_master_rdata),   //               .rdata
		.h2f_RRESP   (axi_master_rresp),   //               .rresp
		.h2f_RLAST   (axi_master_rlast),   //               .rlast
		.h2f_RVALID  (axi_master_rvalid),  //               .rvalid
		.h2f_RREADY  (axi_master_rready)   //               .rready
	);

endmodule
